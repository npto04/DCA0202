library ieee;
use ieee.std_logic_1164.all;

entity cont is
	generic(n : integer := 6);
	port( limite : in std_logic_vector(n-1 downto 0);
			clk : in std_logic;
			saida : out std_logic_vector(n-1 downto 0));
end cont;



architecture arq of cont is
	component reg is
		generic(n : integer := 6);
		port( entrada : in std_logic_vector(n-1 downto 0);
				ld, clk, clr : in std_logic;
				saida : out std_logic_vector(n-1 downto 0));
	end component; 

	component soma is
		generic(n : integer := 4);
		port (		  
				  a,b: in std_logic_vector(n-1 downto 0);
				  s: out std_logic_vector(n-1 downto 0)
			 );
	end component;

	component comp is
		generic(n : integer := 4);
		port (			  
				  a, b: in std_logic_vector(n-1 downto 0);
				  s: out std_logic
			 );
	end component;
	
	signal num1 : std_logic_vector(n-1 downto 0) := (others => '0');
	signal num2 : std_logic_vector(n-1 downto 0);
	signal parar, clr: std_logic;
	signal ld : std_logic := '1';
	signal b : std_logic_vector(n-1 downto 0) := (others => '0');
	
	begin
		b(0) <= '1';
		i1: soma generic map (n) port map (num1,b,num2);
		i2: reg generic map (n) port map(num2,ld,clk,clr,num1);
		i3: comp generic map (n) port map(num1,limite,parar);
		clr <= not parar;
		saida <= num1;
		
end arq;